entity codem_b_l is
   port (
      daytime : in      bit;
      code    : in      bit_vector(3 downto 0);
      reset   : in      bit;
      clk     : in      bit;
      vdd     : in      bit;
      vss     : in      bit;
      door    : out     bit;
      alarm   : out     bit
 );
end codem_b_l;

architecture structural of codem_b_l is
Component nao22_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component a2_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component o4_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component inv_x2
   port (
      i   : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component inv_x8
   port (
      i   : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component o3_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component an12_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component no4_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component sff1_x4
   port (
      ck  : in      bit;
      i   : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component a3_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component na2_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component na3_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component o2_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component on12_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component na4_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      i3  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component oa22_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component no2_x1
   port (
      i0  : in      bit;
      i1  : in      bit;
      nq  : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component ao22_x2
   port (
      i0  : in      bit;
      i1  : in      bit;
      i2  : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

Component buf_x2
   port (
      i   : in      bit;
      q   : out     bit;
      vdd : in      bit;
      vss : in      bit
 );
end component;

signal code_cs           : bit_vector( 2 downto 0);
signal not_code          : bit_vector( 2 downto 1);
signal not_code_cs       : bit_vector( 2 downto 1);
signal on12_x1_sig       : bit;
signal on12_x1_3_sig     : bit;
signal on12_x1_2_sig     : bit;
signal oa22_x2_sig       : bit;
signal o4_x2_sig         : bit;
signal o3_x2_sig         : bit;
signal o2_x2_sig         : bit;
signal o2_x2_3_sig       : bit;
signal o2_x2_2_sig       : bit;
signal not_aux8          : bit;
signal not_aux3          : bit;
signal not_aux2          : bit;
signal not_aux19         : bit;
signal not_aux17         : bit;
signal not_aux11         : bit;
signal not_aux0          : bit;
signal no4_x1_sig        : bit;
signal no2_x1_sig        : bit;
signal no2_x1_3_sig      : bit;
signal no2_x1_2_sig      : bit;
signal na4_x1_sig        : bit;
signal na3_x1_sig        : bit;
signal na3_x1_3_sig      : bit;
signal na3_x1_2_sig      : bit;
signal na2_x1_sig        : bit;
signal na2_x1_2_sig      : bit;
signal mbk_buf_not_aux11 : bit;
signal aux19             : bit;
signal aux18             : bit;
signal aux1              : bit;
signal an12_x1_sig       : bit;
signal a3_x2_sig         : bit;
signal a3_x2_2_sig       : bit;

begin

on12_x1_ins : on12_x1
   port map (
      i0  => code(3),
      i1  => daytime,
      q   => on12_x1_sig,
      vdd => vdd,
      vss => vss
   );

a3_x2_ins : a3_x2
   port map (
      i0  => code(2),
      i1  => not_aux0,
      i2  => on12_x1_sig,
      q   => a3_x2_sig,
      vdd => vdd,
      vss => vss
   );

not_aux8_ins : nao22_x1
   port map (
      i0  => code_cs(2),
      i1  => code(3),
      i2  => a3_x2_sig,
      nq  => not_aux8,
      vdd => vdd,
      vss => vss
   );

not_aux0_ins : a2_x2
   port map (
      i0  => code(0),
      i1  => not_code(1),
      q   => not_aux0,
      vdd => vdd,
      vss => vss
   );

na3_x1_ins : na3_x1
   port map (
      i0  => code(3),
      i1  => not_code(2),
      i2  => aux1,
      nq  => na3_x1_sig,
      vdd => vdd,
      vss => vss
   );

not_aux11_ins : o2_x2
   port map (
      i0  => code_cs(2),
      i1  => na3_x1_sig,
      q   => not_aux11,
      vdd => vdd,
      vss => vss
   );

o4_x2_ins : o4_x2
   port map (
      i0  => code(0),
      i1  => code(1),
      i2  => reset,
      i3  => code(3),
      q   => o4_x2_sig,
      vdd => vdd,
      vss => vss
   );

not_aux17_ins : o4_x2
   port map (
      i0  => o4_x2_sig,
      i1  => code(2),
      i2  => code_cs(2),
      i3  => not_code_cs(1),
      q   => not_aux17,
      vdd => vdd,
      vss => vss
   );

not_code_cs_1_ins : inv_x2
   port map (
      i   => code_cs(1),
      nq  => not_code_cs(1),
      vdd => vdd,
      vss => vss
   );

not_aux19_ins : inv_x2
   port map (
      i   => aux19,
      nq  => not_aux19,
      vdd => vdd,
      vss => vss
   );

not_aux3_ins : o2_x2
   port map (
      i0  => not_aux2,
      i1  => not_code_cs(2),
      q   => not_aux3,
      vdd => vdd,
      vss => vss
   );

not_code_cs_2_ins : inv_x2
   port map (
      i   => code_cs(2),
      nq  => not_code_cs(2),
      vdd => vdd,
      vss => vss
   );

not_aux2_ins : on12_x1
   port map (
      i0  => aux1,
      i1  => code(3),
      q   => not_aux2,
      vdd => vdd,
      vss => vss
   );

not_code_2_ins : inv_x2
   port map (
      i   => code(2),
      nq  => not_code(2),
      vdd => vdd,
      vss => vss
   );

not_code_1_ins : inv_x8
   port map (
      i   => code(1),
      nq  => not_code(1),
      vdd => vdd,
      vss => vss
   );

aux19_ins : no2_x1
   port map (
      i0  => reset,
      i1  => code_cs(0),
      nq  => aux19,
      vdd => vdd,
      vss => vss
   );

aux18_ins : an12_x1
   port map (
      i0  => reset,
      i1  => code_cs(0),
      q   => aux18,
      vdd => vdd,
      vss => vss
   );

aux1_ins : no2_x1
   port map (
      i0  => code(0),
      i1  => not_code(1),
      nq  => aux1,
      vdd => vdd,
      vss => vss
   );

o3_x2_ins : o3_x2
   port map (
      i0  => not_aux19,
      i1  => not_aux3,
      i2  => not_code(2),
      q   => o3_x2_sig,
      vdd => vdd,
      vss => vss
   );

na2_x1_ins : na2_x1
   port map (
      i0  => not_aux17,
      i1  => o3_x2_sig,
      nq  => na2_x1_sig,
      vdd => vdd,
      vss => vss
   );

code_cs_0_ins : sff1_x4
   port map (
      ck  => clk,
      i   => na2_x1_sig,
      q   => code_cs(0),
      vdd => vdd,
      vss => vss
   );

an12_x1_ins : an12_x1
   port map (
      i0  => mbk_buf_not_aux11,
      i1  => aux18,
      q   => an12_x1_sig,
      vdd => vdd,
      vss => vss
   );

code_cs_1_ins : sff1_x4
   port map (
      ck  => clk,
      i   => an12_x1_sig,
      q   => code_cs(1),
      vdd => vdd,
      vss => vss
   );

o2_x2_ins : o2_x2
   port map (
      i0  => code(2),
      i1  => not_aux2,
      q   => o2_x2_sig,
      vdd => vdd,
      vss => vss
   );

no4_x1_ins : no4_x1
   port map (
      i0  => code_cs(1),
      i1  => o2_x2_sig,
      i2  => code_cs(2),
      i3  => not_aux19,
      nq  => no4_x1_sig,
      vdd => vdd,
      vss => vss
   );

on12_x1_2_ins : on12_x1
   port map (
      i0  => not_aux17,
      i1  => no4_x1_sig,
      q   => on12_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

code_cs_2_ins : sff1_x4
   port map (
      ck  => clk,
      i   => on12_x1_2_sig,
      q   => code_cs(2),
      vdd => vdd,
      vss => vss
   );

o2_x2_2_ins : o2_x2
   port map (
      i1  => not_aux11,
      i0  => code_cs(1),
      q   => o2_x2_2_sig,
      vdd => vdd,
      vss => vss
   );

a3_x2_2_ins : a3_x2
   port map (
      i0  => aux18,
      i1  => not_aux8,
      i2  => o2_x2_2_sig,
      q   => a3_x2_2_sig,
      vdd => vdd,
      vss => vss
   );

no2_x1_ins : no2_x1
   port map (
      i0  => code(0),
      i1  => code(3),
      nq  => no2_x1_sig,
      vdd => vdd,
      vss => vss
   );

oa22_x2_ins : oa22_x2
   port map (
      i0  => not_code_cs(2),
      i1  => no2_x1_sig,
      i2  => code(2),
      q   => oa22_x2_sig,
      vdd => vdd,
      vss => vss
   );

no2_x1_2_ins : no2_x1
   port map (
      i0  => code(2),
      i1  => not_code(1),
      nq  => no2_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

na2_x1_2_ins : na2_x1
   port map (
      i0  => no2_x1_2_sig,
      i1  => code_cs(1),
      nq  => na2_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_3_ins : na3_x1
   port map (
      i0  => daytime,
      i1  => code(3),
      i2  => not_aux0,
      nq  => na3_x1_3_sig,
      vdd => vdd,
      vss => vss
   );

na3_x1_2_ins : na3_x1
   port map (
      i0  => code(2),
      i1  => not_aux3,
      i2  => na3_x1_3_sig,
      nq  => na3_x1_2_sig,
      vdd => vdd,
      vss => vss
   );

o2_x2_3_ins : o2_x2
   port map (
      i0  => code(1),
      i1  => code(2),
      q   => o2_x2_3_sig,
      vdd => vdd,
      vss => vss
   );

on12_x1_3_ins : on12_x1
   port map (
      i0  => not_code_cs(1),
      i1  => o2_x2_3_sig,
      q   => on12_x1_3_sig,
      vdd => vdd,
      vss => vss
   );

na4_x1_ins : na4_x1
   port map (
      i0  => on12_x1_3_sig,
      i1  => na3_x1_2_sig,
      i2  => na2_x1_2_sig,
      i3  => oa22_x2_sig,
      nq  => na4_x1_sig,
      vdd => vdd,
      vss => vss
   );

alarm_ins : oa22_x2
   port map (
      i0  => na4_x1_sig,
      i1  => aux19,
      i2  => a3_x2_2_sig,
      q   => alarm,
      vdd => vdd,
      vss => vss
   );

no2_x1_3_ins : no2_x1
   port map (
      i0  => reset,
      i1  => not_aux8,
      nq  => no2_x1_3_sig,
      vdd => vdd,
      vss => vss
   );

door_ins : ao22_x2
   port map (
      i0  => code_cs(0),
      i1  => code(3),
      i2  => no2_x1_3_sig,
      q   => door,
      vdd => vdd,
      vss => vss
   );

mbk_buf_not_aux111 : buf_x2
   port map (
      i   => not_aux11,
      q   => mbk_buf_not_aux11,
      vdd => vdd,
      vss => vss
   );


end structural;
